--=========================================================================================
--
--   ░█▀█░▀█▀░█▀█░█▀█░█▀█░█▀▀░█░░░█▀▀░░░█░█░█░█░░░█▀▀░█▀▄░█▀█░█░█░█▀█░░░░░░░█░░░█░░░█▀▀
--   ░█▀▀░░█░░█░█░█░█░█▀█░█░░░█░░░█▀▀░░░█▀█░█▄█░░░█░█░█▀▄░█░█░█░█░█▀▀░░░░░░░█░░░█░░░█░░
--   ░▀░░░▀▀▀░▀░▀░▀░▀░▀░▀░▀▀▀░▀▀▀░▀▀▀░░░▀░▀░▀░▀░░░▀▀▀░▀░▀░▀▀▀░▀▀▀░▀░░░▄▀░░░░▀▀▀░▀▀▀░▀▀▀
--
--
-- File Name     : my_module.vhd
-- Author        : your name           
-- Project       : project name
-- HDL Version   : version                
-- Description   : brief explanation of what module does 
--                 
-- Dependencies  : List other HDL files, libraries, or packages required
-- Revision      : address to configuration management site
--
--=========================================================================================