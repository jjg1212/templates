--=========================================================================================
--
--   ░█▀█░▀█▀░█▀█░█▀█░█▀█░█▀▀░█░░░█▀▀░░░█░█░█░█░░░█▀▀░█▀▄░█▀█░█░█░█▀█░░░░░░░█░░░█░░░█▀▀
--   ░█▀▀░░█░░█░█░█░█░█▀█░█░░░█░░░█▀▀░░░█▀█░█▄█░░░█░█░█▀▄░█░█░█░█░█▀▀░░░░░░░█░░░█░░░█░░
--   ░▀░░░▀▀▀░▀░▀░▀░▀░▀░▀░▀▀▀░▀▀▀░▀▀▀░░░▀░▀░▀░▀░░░▀▀▀░▀░▀░▀▀▀░▀▀▀░▀░░░▄▀░░░░▀▀▀░▀▀▀░▀▀▀
--
--
-- File Name     : my_module.vhd
-- Author        : your name           
-- Project       : project name
-- HDL Version   : version                
-- Description   : brief explanation of what module does 
--                 
-- Dependencies  : List other HDL files, libraries, or packages required
-- Revision      : address to configuration management site
--
--=========================================================================================

library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;

entity <my_module> is
	   generic(
		   	
		   );
		   port(
			         
			   );
		end <my_module>;
		
		architecture rtl of <my_module> is
			
			
			begin
				
				
			end architecture;